
package reset_pkg is

  type reset_type is (none, sync, async);   

end reset_pkg;
 
  